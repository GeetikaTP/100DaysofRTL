module fulladder_tb();

reg a,b,c;
wire sum,carry;

fulladder uut(a,b,c,sum,carry);

initial begin
#10;
a=1'b0; b=1'b0; c=1'b0;
#10;
a=1'b0; b=1'b0; c=1'b1;
#10;
a=1'b0; b=1'b1; c=1'b0;
#10;
a=1'b0; b=1'b1; c=1'b1;
#10;
a=1'b1; b=1'b0; c=1'b0;
#10;
a=1'b1; b=1'b0; c=1'b1;
#10;
a=1'b1; b=1'b1; c=1'b0;
#10;
a=1'b1; b=1'b1; c=1'b1;
#10;
end
endmodule
